`include "./src/common_usr/avl_stream_if.vh"
`include "./src/struct_s.sv"

// nf submodule
module bypass_front_avlstrm (
    input logic Clk, 
    input logic Rst_n,

    avl_stream_if.rx in_pkt,
    avl_stream_if.rx in_meta,
    avl_stream_if.rx in_usr,
    avl_stream_if.tx out_pkt,
    avl_stream_if.tx out_meta,
    avl_stream_if.tx out_usr,
    avl_stream_if.tx bypass_pkt,
    avl_stream_if.tx bypass_meta,
    avl_stream_if.tx bypass_usr
);

bypass_nf_front bypass_nf_front_inst(
    .clk                    (Clk),
    .rst                    (~Rst_n),
    .in_pkt_sop             (in_pkt.sop),
    .in_pkt_eop             (in_pkt.eop),
    .in_pkt_data            (in_pkt.data),
    .in_pkt_empty           (in_pkt.empty),
    .in_pkt_valid           (in_pkt.valid),
    .in_pkt_ready           (in_pkt.ready),
    .in_pkt_almost_full     (),
    .in_meta_valid          (in_meta.valid),
    .in_meta_ready          (in_meta.ready),
    .in_meta_data           (in_meta.data),
    .in_meta_almost_full    (),
    .in_usr_sop             (in_usr.sop),
    .in_usr_eop             (in_usr.eop),
    .in_usr_data            (in_usr.data),
    .in_usr_empty           (in_usr.empty),
    .in_usr_valid           (in_usr.valid),
    .in_usr_ready           (in_usr.ready),
    .in_usr_almost_full     (),
    .out_pkt_data           (out_pkt.data),
    .out_pkt_sop            (out_pkt.sop),
    .out_pkt_eop            (out_pkt.eop),
    .out_pkt_empty          (out_pkt.empty),
    .out_pkt_valid          (out_pkt.valid),
    .out_pkt_ready          (out_pkt.ready),
    .out_pkt_almost_full    (out_pkt.almost_full),
    .out_pkt_channel        (out_pkt.channel),
    .out_meta_data          (out_meta.data),
    .out_meta_valid         (out_meta.valid),
    .out_meta_ready         (out_meta.ready),
    .out_meta_almost_full   (out_meta.almost_full),
    .out_meta_channel       (),
    .out_usr_data           (out_usr.data),
    .out_usr_sop            (out_usr.sop),
    .out_usr_eop            (out_usr.eop),
    .out_usr_empty          (out_usr.empty),
    .out_usr_valid          (out_usr.valid),
    .out_usr_ready          (out_usr.ready),
    .out_usr_almost_full    (out_usr.almost_full),
    .out_usr_channel        (),
    .bypass_pkt_data           (bypass_pkt.data),
    .bypass_pkt_sop            (bypass_pkt.sop),
    .bypass_pkt_eop            (bypass_pkt.eop),
    .bypass_pkt_empty          (bypass_pkt.empty),
    .bypass_pkt_valid          (bypass_pkt.valid),
    .bypass_pkt_ready          (bypass_pkt.ready),
    .bypass_pkt_almost_full    (bypass_pkt.almost_full),
    .bypass_pkt_channel        (),
    .bypass_meta_data          (bypass_meta.data),
    .bypass_meta_valid         (bypass_meta.valid),
    .bypass_meta_ready         (bypass_meta.ready),
    .bypass_meta_almost_full   (bypass_meta.almost_full),
    .bypass_meta_channel       (),
    .bypass_usr_data           (bypass_usr.data),
    .bypass_usr_sop            (bypass_usr.sop),
    .bypass_usr_eop            (bypass_usr.eop),
    .bypass_usr_empty          (bypass_usr.empty),
    .bypass_usr_valid          (bypass_usr.valid),
    .bypass_usr_ready          (bypass_usr.ready),
    .bypass_usr_almost_full    (bypass_usr.almost_full),
    .bypass_usr_channel        ()
);

endmodule

module bypass_front_avlstrm_round_robin (
    input logic Clk, 
    input logic Rst_n,

    avl_stream_if.rx in_pkt,
    avl_stream_if.rx in_meta,
    avl_stream_if.rx in_usr,
    avl_stream_if.tx out_pkt,
    avl_stream_if.tx out_meta,
    avl_stream_if.tx out_usr,
    avl_stream_if.tx bypass_pkt,
    avl_stream_if.tx bypass_meta,
    avl_stream_if.tx bypass_usr
);

bypass_nf_front_rr bypass_nf_front_inst(
    .clk                    (Clk),
    .rst                    (~Rst_n),
    .in_pkt_sop             (in_pkt.sop),
    .in_pkt_eop             (in_pkt.eop),
    .in_pkt_data            (in_pkt.data),
    .in_pkt_empty           (in_pkt.empty),
    .in_pkt_valid           (in_pkt.valid),
    .in_pkt_ready           (in_pkt.ready),
    .in_pkt_almost_full     (),
    .in_meta_valid          (in_meta.valid),
    .in_meta_ready          (in_meta.ready),
    .in_meta_data           (in_meta.data),
    .in_meta_almost_full    (),
    .in_usr_sop             (in_usr.sop),
    .in_usr_eop             (in_usr.eop),
    .in_usr_data            (in_usr.data),
    .in_usr_empty           (in_usr.empty),
    .in_usr_valid           (in_usr.valid),
    .in_usr_ready           (in_usr.ready),
    .in_usr_almost_full     (),
    .out_pkt_data           (out_pkt.data),
    .out_pkt_sop            (out_pkt.sop),
    .out_pkt_eop            (out_pkt.eop),
    .out_pkt_empty          (out_pkt.empty),
    .out_pkt_valid          (out_pkt.valid),
    .out_pkt_ready          (out_pkt.ready),
    .out_pkt_almost_full    (out_pkt.almost_full),
    .out_pkt_channel        (out_pkt.channel),
    .out_meta_data          (out_meta.data),
    .out_meta_valid         (out_meta.valid),
    .out_meta_ready         (out_meta.ready),
    .out_meta_almost_full   (out_meta.almost_full),
    .out_meta_channel       (),
    .out_usr_data           (out_usr.data),
    .out_usr_sop            (out_usr.sop),
    .out_usr_eop            (out_usr.eop),
    .out_usr_empty          (out_usr.empty),
    .out_usr_valid          (out_usr.valid),
    .out_usr_ready          (out_usr.ready),
    .out_usr_almost_full    (out_usr.almost_full),
    .out_usr_channel        (),
    .bypass_pkt_data           (bypass_pkt.data),
    .bypass_pkt_sop            (bypass_pkt.sop),
    .bypass_pkt_eop            (bypass_pkt.eop),
    .bypass_pkt_empty          (bypass_pkt.empty),
    .bypass_pkt_valid          (bypass_pkt.valid),
    .bypass_pkt_ready          (bypass_pkt.ready),
    .bypass_pkt_almost_full    (bypass_pkt.almost_full),
    .bypass_pkt_channel        (),
    .bypass_meta_data          (bypass_meta.data),
    .bypass_meta_valid         (bypass_meta.valid),
    .bypass_meta_ready         (bypass_meta.ready),
    .bypass_meta_almost_full   (bypass_meta.almost_full),
    .bypass_meta_channel       (),
    .bypass_usr_data           (bypass_usr.data),
    .bypass_usr_sop            (bypass_usr.sop),
    .bypass_usr_eop            (bypass_usr.eop),
    .bypass_usr_empty          (bypass_usr.empty),
    .bypass_usr_valid          (bypass_usr.valid),
    .bypass_usr_ready          (bypass_usr.ready),
    .bypass_usr_almost_full    (bypass_usr.almost_full),
    .bypass_usr_channel        ()
);

endmodule
